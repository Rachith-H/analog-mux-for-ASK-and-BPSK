magic
tech scmos
timestamp 1760677986
<< nwell >>
rect -6 18 10 28
rect -6 -20 10 -10
<< polysilicon >>
rect 1 42 3 45
rect 1 36 3 38
rect 1 27 3 29
rect 1 13 3 19
rect 1 4 3 9
rect 1 -2 3 0
rect 1 -11 3 -9
rect 1 -23 3 -19
<< ndiffusion >>
rect -1 38 1 42
rect 3 38 5 42
rect -1 0 1 4
rect 3 0 5 4
<< pdiffusion >>
rect -1 23 1 27
rect -5 19 1 23
rect 3 23 5 27
rect 3 19 9 23
rect -1 -15 1 -11
rect -5 -19 1 -15
rect 3 -15 5 -11
rect 3 -19 9 -15
<< metal1 >>
rect -4 45 -1 49
rect -5 35 -1 38
rect -10 31 -1 35
rect -5 27 -1 31
rect 5 35 9 38
rect 5 31 17 35
rect 5 27 9 31
rect 13 13 17 31
rect -7 9 -1 13
rect 13 9 21 13
rect -5 -3 -1 0
rect -10 -7 -1 -3
rect -5 -11 -1 -7
rect 5 -3 9 0
rect 13 -3 17 9
rect 5 -7 17 -3
rect 5 -11 9 -7
rect -4 -27 -1 -23
<< ntransistor >>
rect 1 38 3 42
rect 1 0 3 4
<< ptransistor >>
rect 1 19 3 27
rect 1 -19 3 -11
<< polycontact >>
rect -1 45 3 49
rect -1 9 3 13
rect -1 -27 3 -23
<< ndcontact >>
rect -5 38 -1 42
rect 5 38 9 42
rect -5 0 -1 4
rect 5 0 9 4
<< pdcontact >>
rect -5 23 -1 27
rect 5 23 9 27
rect -5 -15 -1 -11
rect 5 -15 9 -11
<< labels >>
rlabel metal1 -10 31 -10 35 3 in1
rlabel metal1 -10 -7 -10 -3 3 in2
rlabel metal1 -7 9 -7 13 3 selbar
rlabel metal1 -4 -27 -4 -23 1 sel
rlabel metal1 -4 45 -4 49 1 sel
rlabel metal1 21 9 21 13 7 out
<< end >>
